// `include "defines.v"

// ID 模块的作用是对指令进行译码，得到最终运算的类型、子类型、源操作数1、源操作数2、要写入的目的寄存器地址等信息
// 运算类型：逻辑运算、移位运算、算术运算等
// 子类型： 更加详细的运算类型。比如: 当运算类型是逻辑运算时，运算子类型可以是逻辑“或”、逻辑“与”、逻辑“异或”运算
module id(

	input wire  rst,                        // 复位信号
	input wire[`InstAddrBus]    pc_i,       // 译码阶段的指令对应的地址
	input wire[`InstBus]    inst_i,         // 译码阶段的指令

	input wire[`RegBus] reg1_data_i,        // 从Regfile输入的第一个读寄存器端口的输入
	input wire[`RegBus] reg2_data_i,        // 从Regfile输入的第二个读寄存器端口的输入

	//送到regfile的信息
	output reg  reg1_read_o,                // Regfile模块的第一个读寄存器端口的读使能信号
	output reg  reg2_read_o,                // Regfile模块的第二个读寄存器端口的读使能信号
	output reg[`RegAddrBus] reg1_addr_o,    // Regfile模块的第一个读寄存器端口的读地址信号
	output reg[`RegAddrBus] reg2_addr_o, 	// Regfile模块的第二个读寄存器端口的读地址信号     
	
	//送到执行阶段的信息
	output reg[`AluOpBus]   aluop_o,        // 译码阶段的指令要进行的运算的子类型
	output reg[`AluSelBus]  alusel_o,       // 译码阶段的指令要进行的运算的类型   
	output reg[`RegBus] reg1_o,             // 译码阶段的指令要进行的运算的源操作数1
	output reg[`RegBus] reg2_o,             // 译码阶段的指令要进行的运算的源操作数2
	output reg[`RegAddrBus] wd_o,           // 译码阶段的指令要写入的目的寄存器地址
	output reg  wreg_o                      // 译码阶段的指令是否有要写入的目的寄存器
);

    // 取得指令的指令码，功能吗
    // 对于ori只需要通过判断第26-31bit的值，即可判断是否是ori指令
    wire[5:0] op = inst_i[31:26];
    wire[4:0] op2 = inst_i[10:6];
    wire[5:0] op3 = inst_i[5:0];
    wire[4:0] op4 = inst_i[20:16];

    // 保存指令执行需要的立即数
    reg[`RegBus]	imm;
    // 指示指令是否有效
    reg instvalid;
  
    // 第一阶段: 对指令进行译码。依据指令中的特征字段区分指令，对指令ori而言，只需要识别26-31bit的指令码是否为6'b001101
    // 即可判断是否是ori指令，其中的宏定义EXE_ORI就是6‘b001101,op就是指令的26-31bit
    // 所以当op等于EXE_ORI时，就表示是ori指令
	always @ (*) begin	
		if (rst == `RstEnable) begin
			aluop_o <= `EXE_NOP_OP;
			alusel_o <= `EXE_RES_NOP;
			wd_o <= `NOPRegAddr;
			wreg_o <= `WriteDisable;
			instvalid <= `InstValid;
			reg1_read_o <= 1'b0;
			reg2_read_o <= 1'b0;
			reg1_addr_o <= `NOPRegAddr;
			reg2_addr_o <= `NOPRegAddr;
			imm <= 32'h0;			
	  	end else begin
			aluop_o <= `EXE_NOP_OP;
			alusel_o <= `EXE_RES_NOP;
			wd_o <= inst_i[15:11];
			wreg_o <= `WriteDisable;
			instvalid <= `InstInvalid;	   
			reg1_read_o <= 1'b0;
			reg2_read_o <= 1'b0;
			reg1_addr_o <= inst_i[25:21];   //默认通过Regfile读端口1读取的寄存器地址
			reg2_addr_o <= inst_i[20:16];	//默认通过Regfile读端口2读取的寄存器地址
			imm <= `ZeroWord;

            case (op)
                `EXE_ORI: begin   // ORI指令。根据op的值判断是否是ori指令
                    // ori指令需要将结果写入目的寄存器，所以wreg_o为WriteEnable
                    wreg_o <= `WriteEnable;
                    // 运算的子类型是逻辑“或”运算
                    aluop_o <= `EXE_OR_OP;
                    // 运算类型是逻辑运算
                    alusel_o <= `EXE_RES_LOGIC; 
                    // 需要通过Regfile的读端口1读取寄存器
                    reg1_read_o <= 1'b1;
                    // 不需要通过Regfile的读端口2读取寄存器
                    reg2_read_o <= 1'b0;
                    // 指令执行需要的立即数
                    imm <= {16'h0, inst_i[15:0]};
                    // 指令执行要写的目睹寄存器地址
                    wd_o <= inst_i[20:16];
                    // ori指令是有效指令
                    instvalid <= `InstValid;	
                end 							 
                default: begin
                end
            endcase		  // case op			
		end       // if
	end         // always
	

    // 第二阶段: 确定进行运算的源操作数1
    // 如果reg1_read_o为1，那么就将从Regfile模块读端口1读取的寄存器的值作为源操作数1
    // 如果reg1_read_o 为0，那么久将立即数作为源操作数1，对于ori而言，此处选择从Regfile模块读端口1读取的寄存器的值作为源操作数1
    // 该值将通过reg1_o 端口被传递到执行阶段
	always @ (*) begin
		if(rst == `RstEnable) begin
			reg1_o <= `ZeroWord;
	    end else if(reg1_read_o == 1'b1) begin
	  	    reg1_o <= reg1_data_i;  // Regfile 读端口1的输出值
	    end else if(reg1_read_o == 1'b0) begin
	  	    reg1_o <= imm;  // 立即数
	    end else begin
	        reg1_o <= `ZeroWord;
	  end
	end
    
    // 第三阶段: 确定进行运算的源操作数2
    // 如果reg2_read_o为1，那么就将从Regfile模块读端口2读取的寄存器的值作为源操作数2
    // 如果reg2_read_o 为0，那么久将立即数作为源操作数2，对于ori而言，此处选择从Regfile模块读端口1读取的寄存器的值作为源操作数2
    // 该值将通过reg2_o 端口被传递到执行阶段
	always @ (*) begin
		if(rst == `RstEnable) begin
			reg2_o <= `ZeroWord;
	    end else if(reg2_read_o == 1'b1) begin
	  	    reg2_o <= reg2_data_i;  // Regfile 读端口2的输出值
	    end else if(reg2_read_o == 1'b0) begin
	  	    reg2_o <= imm;          // 立即数
	    end else begin
	        reg2_o <= `ZeroWord;
	    end
	end

endmodule